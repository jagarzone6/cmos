* Simulación Circuito Del ejercicio 5.5-20 Allen CMOS Amplifier Class A
* Usando modelo de canal largo y modelo simple, con parametros del allen
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A
////////////------////////////////////

*Circuito A modelo que incluye lamba, nivel 3 canal largo
*vout
VDD VDD 0 DC 2 AC 0
Vss Vss 0 DC -2 AC 0
Vgg2 gateM2 0 DC 0 AC 0

M2 out gateM2 vdd VDD pmoslevel3 W=13609u L=1u
M1 out vin vss Vss nmoslevel3 W=5971u L=1u

*Resistor de carga y capacitor de carga
Rl out 0 100
Cl out 0 1n


*///Voltaje de entrada vin AC y DC para ambos circuitos/////
* Voltaje DC de vin
VGin VGcommon11 0 DC 0 AC 0
*Fuente AC en los gates despues de la fuente DC de polarizacion
VO vin VGcommon11 sin(0 1 10k) dc=0 ac=1


.model nmoslevel3 nmos LEVEL=3
+ Vto=0.5 KP=100E-6 gamma=0.5 phi=0.7
+ DELTA=3.0 U0=650 ETA=3E-6 KAPPA=0.3 THETA=0.1
+ TOX=200E-10 NSUB=1E17 XJ=500E-9 LD=100E-9 NFS=1E12
+ cgso=200E-12 cgdo=200E-12 cgbo=1E-10
+ cj=400E-6 cjsw=300E-12 mj=0.5 mjsw=0.5
+ RSH=0 VMAX=1E5 TPG=1 PB=1

.model pmoslevel3 pmos LEVEL=3
+ Vto=-0.5 KP=50E-6 gamma=0.6 phi=0.7
+ DELTA=0.1 U0=250 ETA=0 KAPPA=1 THETA=0.1
+ TOX=200E-10 NSUB=1E17 XJ=500E-9 LD=100E-9 NFS=1E12
+ cgso=200E-12 cgdo=200E-12 cgbo=1E-10
+ cj=400E-6 cjsw=300E-12 mj=0.5 mjsw=0.5
+ RSH=0 VMAX=5E4 TPG=1 PB=1


.control
set color0 =white
set color1=black
op
show all

*Ganacia en AC barrido en frecuencia vout/vin AC
ac dec 10 1 10ghz
*Ganancia en decibeles
plot db(mag(v(out))/mag(v(vgcommon11,vin)))
*Ganancia en magnitud V/V
plot mag(v(out))/mag(v(vgcommon11,vin))

*Transitorio
tran .000001s .001s

*Corrientes de polarizacion DC del transistor M2
plot i(vdd)

*Voltaje de entrada AC v(vgcommon112,vin2)
plot v(vgcommon11,vin)
*voltaje de salida AC v(out)
plot v(out)



.endc