* Simulación Circuito De las figuras 4,1,12_13 CMOS Switch Level 1
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

VDD VDD 0 DC 5 AC 0
Vin Vin 0 DC 3 AC 0
RL RLo 0 0.00000001
VRL SOURCE RLo DC 0 AC 0
M1 Vin VDD SOURCE 0 nmoslevel1 W=60 L=2
M2 Vin 0 SOURCE 0 pmoslevel1 W=60 L=2


.model nmoslevel1 nmos LEVEL=1 Vto=0.8 KP=120u LAMBDA=0.01 U0=650
.model pmoslevel1 pmos LEVEL=1 Vto=-0.9 KP=40u LAMBDA=0.0125 U0=250

.control
set color0 =white
set color1=black
op
show all
dc vin 0 5 0.01
plot vin/i(vrl)
.endc
