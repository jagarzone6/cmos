*** SPICE deck for cell Current_mirror_bias_SIM{sch} from library Fig-20-25-Sim
*** Created on Mon Oct 03, 2016 12:52:34
*** Last revised on Mon Oct 03, 2016 13:58:16
*** Written on Mon Oct 03, 2016 13:58:31 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
*.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
*+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
*+LVLCOD=1
.MODEL Nmodel NMOS LEVEL=3
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL Pmodel PMOS LEVEL=3
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd
*** WARNING: no power connection for P-transistor wells in cell 'Current_mirror_bias_SIM{sch}'

*** TOP LEVEL CELL: Current_mirror_bias_SIM{sch}

* Spice Declaration nodes in cell cell 'Current_mirror_bias_SIM{sch}'
Vdd VDDin gnd 5
.dc Vdd 0 6 1m
.include long_channel_3_models.txt
Mnmos@0 gnd net@0 net@2 gnd Nmodel L=2U W=10U
Mnmos@1 gnd net@0 net@0 gnd Nmodel L=2U W=10U
Mnmos@2 net@9 net@2 net@0 gnd Nmodel L=1U W=10U
Mnmos@3 net@9 net@0 net@20 gnd Nmodel L=2U W=40U
Mpmos@0 net@2 net@2 net@8 VDDin Pmodel L=100U W=10U
Mpmos@1 net@0 net@9 net@8 VDDin Pmodel L=2U W=30U
Mpmos@2 net@8 net@9 net@9 VDDin Pmodel L=2U W=30U
Rres@0 net@20 gnd 6.5k
.END
