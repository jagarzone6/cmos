
* Simulación Circito Número 4 (Espejo de Corriente con Cmos)
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

VDD VDD 0 DC 10 AC 0
VG GATE 0 DC 4 AC 0
RD VDD DRAIN 3000
M1 DRAIN GATE SOURCE 0 nmos W=6 L=2
I1 SOURCE 0 DC 0.002 AC 0
M2 DRAIN2 GATE SOURCE2 0 nmos2 W=6 L=2
I2 SOURCE2 0 DC 0.001 AC 0
.model nmos nmos LEVEL=1 Vto=0.75 KP=120u LAMBDA=0.01 U0=650
.model nmos2 nmos LEVEL=1 Vto=0.75 KP=120u LAMBDA=0.01 U0=650

.control
set color0 =white
set color1=black
op
show all
dc vg 0 5 0.1
plot v(source)
.endc
