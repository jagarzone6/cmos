* Simulación Circuito Espejo de Corriente con Ncmos, valores reales de Kp_n y Vt
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

VDD VDD 0 DC -10 AC 0
V2 VR 0 DC -10 AC 0
VRD RDN VR DC 0 AC 0
RD RDN DRAIN 1000
RP VDD GATE 2000
M1 DRAIN GATE 0 0 pmosideal W=60 L=2
M2 GATE GATE 0 0 pmosideal W=60 L=2

VRD2 RDN2 VR DC 0 AC 0
RD2 RDN2 DRAIN2 1000
RP2 VDD GATE2 2000
M3 DRAIN2 GATE2 0 0 pmos1 W=60 L=2
M4 GATE2 GATE2 0 0 pmos2 W=60 L=2

.model pmosideal pmos LEVEL=1 Vto=-0.9 KP=40u LAMBDA=0.0125 U0=250
.model pmos1 pmos LEVEL=1 Vto=-1.01696 KP=40u LAMBDA=0.0125 U0=250
.model pmos2 pmos LEVEL=1 Vto=-0.98784 KP=40u LAMBDA=0.0125 U0=250

.control
set color0 =white
set color1=black
op
show all
dc vdd -0.8 -12 -0.01
plot i(vrd) i(vrd2)
.endc
