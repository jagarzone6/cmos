* Bogotá 5 de octubre de 2016
* Universidad Nacional de Colombia 
* CMOS Analógico
* Simulación circuito figura 20.14 Baker (pg 624)
* Grupo Jorge Garzón, Esteban Iafrancesco


** PARA LAMBDA=0.01*******************************************************
VDD VDD 0 DC 5 AC 0
*Vbiasp G4 0 
*Vbiasn G2 0
M1 G2 G2 S1 0 nmos W=10 L=2
M2 D2 G2 S1 0 nmos W=10 L=2
M3 G2 G4 VDD VDD pmos W=30 L=2
M4 G4 G4 VDD VDD pmos W=30 L=2
R S7 0 6500

.MODEL NMOS NMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.01 
+ TOX =200E-10
+ PHI =0.7 VTO = 0.8
+ UO = 650 ETA = 3.0E-6
+ KP=120E-6 VMAX =1E5
+ RSH = 0 NFS =1E12
+ XJ = 500E-9LD = 100E-9
+ CGDO =200E-12 CGSO =200E-12 PB = 1
+ CJ = 400E-6
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.5 DELTA = 3.0 THETA = 0.1 KAPPA =0.3
+ TPG = 1 CGBO =1E-10 MJ = 0.5
*
.MODEL PMOS PMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.01 
+ TOX =200E-10
+ PHI = 0.7 VTO = -0.9 ETA = 0
+ UO = 250 VMAX =5E4
+ KP = 40E-6
+ RSH = 0 NFS =1E12 LD = 100E-9
+ XJ = 500E-9 CGSO =200E-12
+ CGDO =200E-12
+ CJ = 400E-6 PB=1
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.6 DELTA =0.1 THETA = 0.1 KAPPA = 1
+ TPG = -1 CGBO =1E-10 MJ = 0.5


.control
set color0 =white
set color1=black
op
show all
dc VDD 0 6 0.2
plot v(G4) v(G2) 
.endc

** PARA LAMBDA=0.1*********************************************************
.MODEL NMOS NMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.1 
+ TOX =200E-10
+ PHI =0.7 VTO = 0.8
+ UO = 650 ETA = 3.0E-6
+ KP=120E-6 VMAX =1E5
+ RSH = 0 NFS =1E12
+ XJ = 500E-9LD = 100E-9
+ CGDO =200E-12 CGSO =200E-12 PB = 1
+ CJ = 400E-6
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.5 DELTA = 3.0 THETA = 0.1 KAPPA =0.3
+ TPG = 1 CGBO =1E-10 MJ = 0.5
*
.MODEL PMOS PMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.01 
+ TOX =200E-10
+ PHI = 0.7 VTO = -0.9 ETA = 0
+ UO = 250 VMAX =5E4
+ KP = 40E-6
+ RSH = 0 NFS =1E12 LD = 100E-9
+ XJ = 500E-9 CGSO =200E-12
+ CGDO =200E-12
+ CJ = 400E-6 PB=1
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.6 DELTA =0.1 THETA = 0.1 KAPPA = 1
+ TPG = -1 CGBO =1E-10 MJ = 0.5


.control
set color0 =white
set color1=black
op
show all
dc VDD 0 6 0.2
plot v(G4) v(G2) 
.endc

** PARA LAMBDA=0.5*********************************************************
.MODEL NMOS NMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.5 
+ TOX =200E-10
+ PHI =0.7 VTO = 0.8
+ UO = 650 ETA = 3.0E-6
+ KP=120E-6 VMAX =1E5
+ RSH = 0 NFS =1E12
+ XJ = 500E-9LD = 100E-9
+ CGDO =200E-12 CGSO =200E-12 PB = 1
+ CJ = 400E-6
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.5 DELTA = 3.0 THETA = 0.1 KAPPA =0.3
+ TPG = 1 CGBO =1E-10 MJ = 0.5
*
.MODEL PMOS PMOS LEVEL = 3 NSUB =1E17 LAMBDA=0.5 
+ TOX =200E-10
+ PHI = 0.7 VTO = -0.9 ETA = 0
+ UO = 250 VMAX =5E4
+ KP = 40E-6
+ RSH = 0 NFS =1E12 LD = 100E-9
+ XJ = 500E-9 CGSO =200E-12
+ CGDO =200E-12
+ CJ = 400E-6 PB=1
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.6 DELTA =0.1 THETA = 0.1 KAPPA = 1
+ TPG = -1 CGBO =1E-10 MJ = 0.5


.control
set color0 =white
set color1=black
op
show all
dc VDD 0 6 0.2
plot v(G4) v(G2) 
.endc
	

