* Simulación Circuito De las figura 5.2-6 Allen CMOS differential amplifier using a current-mirror load
* Usando valores del ejemplo 5.2-2
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

*Definicion del circuito Amplificador diferencial en modo diferencial
*El bulk de M1 y M2 se conecta al source en ves de a vss
VDD VDD 0 DC 2.5 AC 0
VSS VSS 0 DC -2.5 AC 0
M3 gateM3 gateM3 VDD VDD pmoslevel3 W=8u L=1u
M4 drainM4 gateM3 VDD VDD pmoslevel3 W=8u L=1u
M1 gateM3 VGcommon1 sM1 sM1 nmoslevel3 W=40u L=1u
M2 drainM4 VGcommon2 sM2 sM2 nmoslevel3 W=40u L=1u
M5 drainM5 gateM5 iss VSS nmoslevel3 W=82u L=1u

*Iref para la fuente de corriente de 100u Amps
Ro vdd gateM5 43k
M7 gateM5 gateM5 isc VSS nmoslevel3 W=82u L=1u

*Fuentes de voltage de 0v para medir corriente en los tranisitores M7 (Espejo) M1 y M2
VIcs isc VSS DC 0 AC 0
Vrefm2 sM2 drainM5 DC 0 AC 0
Vrefm1 sM1 drainM5 DC 0 AC 0

* Fuente dc 0 volts para medir la corriente Iss en el transistor M5
VIss iss VSS DC 0 AC 0

* Voltaje DC de gateM2 y gateM1
VGcm1 VGcommon11 0 DC 1 AC 0
VGcm2 VGcommon2 0 DC 1 AC 0

*Fuente AC en los gates despues de la fuente DC de polarizacion
VO VGcommon1 VGcommon11 sin(0 0.002 100k) dc=0 ac=0.002

*Capacitor de salida
C2 drainM4 0 5p

.model nmoslevel3 nmos LEVEL=3
+ Vto=0.8 KP=120E-6 gamma=0.5 phi=0.7
+ DELTA=3.0 U0=650 ETA=3E-6 KAPPA=0.3 THETA=0.1
+ TOX=200E-10 NSUB=1E17 XJ=500E-9 LD=100E-9 NFS=1E12
+ cgso=200E-12 cgdo=200E-12 cgbo=1E-10
+ cj=400E-6 cjsw=300E-12 mj=0.5 mjsw=0.5
+ RSH=0 VMAX=1E5 TPG=1 PB=1

.model pmoslevel3 pmos LEVEL=3
+ Vto=-0.9 KP=40E-6 gamma=0.6 phi=0.7
+ DELTA=0.1 U0=250 ETA=0 KAPPA=1 THETA=0.1
+ TOX=200E-10 NSUB=1E17 XJ=500E-9 LD=100E-9 NFS=1E12
+ cgso=200E-12 cgdo=200E-12 cgbo=1E-10
+ cj=400E-6 cjsw=300E-12 mj=0.5 mjsw=0.5
+ RSH=0 VMAX=5E4 TPG=1 PB=1

.control
set color0 =white
set color1=black
op
show all

*Ganacia en AC barrido en frecuencia vout/vin AC
ac dec 10 1 0.1ghz
plot db(mag(v(drainm4))/mag(v(vgcommon11,vgcommon1)))

*Transitorio
tran .0000001s .0001s

*Corrientes de polarizacion Iss y Idm2 Idm1
plot i(viss) i(vrefm1) i(vrefm2)

*Voltaje de entrada
plot v(vgcommon11,vgcommon1)

*voltaje de salida
plot v(drainm4)
.endc