
* Simulación Circito Número 1 (Carga pasiva RL)
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A
* RD = Resistencia de drenador
* RL = Resistencia de Carga
* VO = tension en la carga (RL)


VDD VDD 0 DC 10 AC 0
VG GATE 0 DC 4.0833 AC 0
VO DRAIN 0 DC 8 AC 0
RL DRAIN 0 2000
RD VDD DRAIN 1000
M1 DRAIN GATE SOURCE 0 nmos W=6 L=2
I1 SOURCE 0 DC 0.002 AC 0

.model nmos nmos LEVEL=1 Vto=0.75 KP=120u LAMBDA=0.01 U0=650

.control
OP
show all
DC VG 0 5 0.1
plot V(SOURCE)
.endc
	







