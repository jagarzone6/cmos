* Bogotá 5 de octubre de 2016
* Universidad Nacional de Colombia
* CMOS Analógico
* Simulación circuito figura 20.28 Baker. Espejo de corriente
* Grupo Jorge Garzón, Esteban Iafrancesco

VDD VDD 0 DC 1 AC 0
VO vo 0 sin(0 0.02 5k) dc=0 ac=0.02
MSU2 VDD D1 D1 VDD pmos W=10 L=20
M2 D1 D4 0 0 nmos W=50 L=2
MSU3 G4 D1 D4 0 nmos W=10 L=1
M4 VDD G4 D4 VDD pmos W=100 L=2
M5 D4 D4 0 0 nmos W=50 L=2
M6 VDD G6 G6 VDD pmos W=100 L=2
M7 G6 G7 0 0 nmos W=50 L=2
M8 VDD G6 G4 VDD pmos W=100 L=2
M9 G4 D4 0 0 nmos W=50 L=2
M10 VDD G4 G7 VDD pmos W=100 L=2
M11 G7 G7 S11 0 nmos W=200 L=2
Vrl S11 S12 DC 0 AC 0
Rl S12 0 5500

*Cacodo con una resistencia de 100 ohmios en serie
Roo vo Dcasc 100
MCasc Dcasc D4 Scasc 0 nmos W=50 L=2
VCasc Scasc 0 DC 0 AC 0
*MCasc vo D4 Scasc 0 nmos W=50 L=2
*VCasc Scasc 0 DC 0 AC 0


.MODEL NMOS NMOS   LEVEL   = 54
+binunit = 1 paramchk= 1 mobmod = 0
+capmod = 2 igcmod = 1 igbmod = 1 geomod = 1
+diomod = 1 rdsmod = 0 rbodymod= 1 rgatemod= 1
+permod = 1
+tnom = 27
+epsrox = 3.9
+LL =0
+lw =0
+lwl = 0
+vth0 = 0.22
+k3b = 0
+dvt2 = -0.032
+dsub = 2
+dvtp1 = 0.05
+ngate = 5e+020
+cdsc = 0.0002
+voff =-0.15
+vfb = -0.55
+uc =-3e-011
+a1 =0
+keta = 0.04
+pdiblc1 = 0.028
+pvag = 1e-020
+fprout =0.2
+rsh = 3
+rdswmin = 0
+prwb = 6.8e-011
+beta0 =30
+egidl =0.8
+aigbacc = 0.012
+nigbacc = 1
+eigbinv= 1.1
+cigc = 0.002
+nigc = 1
+xrcrg1 = 12
+cgso =6.238e-010
+cgsl = 2.495e-10
+moin = 15
+kt1 = -0.21
+ua1 = 1e-009
+at = 53000
+fnoimod = 1
+jss = 0.0001
+ijthsfwd= 0.01
+jsd = 0.0001
+ijthdfwd= 0.01
+pbs =1
+cjsws =5e-010
+mjswgs = 0.33
+pbswd = 1
+cjswgd = 5e-010
+tpbsw =0.005
+xtis = 3
+acnqsmod= 0
+toxe = 1.4e-009
+wint = 5e-009
+wl =0
+ww =0
+wwl = 0
+k1 = 0.35
+w0 = 2.5e-006
+dvt0w = 0
+minv = 0.05
+lpe0 = 5.75e-008
+ndep =2.8e+018
+cdscb = 0
+nfactor = 1.2
+u0 = 0.032
+vsat =1.1e+005
+a2 =1
+dwg = 0
+pdiblc2 = 0.022
+delta =0.01
+pdits = 0.2
+rdsw = 150
+rdwmin = 0
+wr =1
+agidl =0.0002
+bigbacc = 0.0028
+aigbinv = 0.014
+nigbinv = 3
+aigsd =0.017
+poxedge = 1
+xrcrg2 = 5
+trnqsmod= 0
+toxp =7e-010
+lint = 1.2e-008
+lln =1
+lwn = 1
+xpart = 0
+k2 = 0.05
+dvt0 = 2.8
+dvt1w =0
+voffl =0
+lpeb =2.3e-010
+nsd =1e+020
+cdscd = 0
+eta0 =0.15
+ua =1.6e-010
+a0 =2
+b0 =-1e-020
+dwb =0
+pdiblcb = -0.005
+pscbe1 = 8.14e+8
+pditsd =0.23
+rsw = 150
+rswmin = 0
+alpha0 =0.074
+bgidl =2.1e+009
+cigbacc = 0.002
+bigbinv = 0.004
+aigc =0.017
+bigsd =0.0028
+pigcd = 1
+cgdo =6.238e-010 cgbo =2.56e-011
+ckappas = 0.02
+noff = 0.9
+kt1l =0.0
+ub1 =-3.5e-019
+tnoimod = 0
+jsws =1e-011
+ijthsrev= 0.001
+jswd =1e-011
+ijthdrev= 0.001
+cjs = 0.0005
+mjsws = 0.33
+pbd =1
+cjswd =5e-010
+mjswgd = 0.33
+tcjsw = 0.001
+xtid = 3
+ckappad = 0.02
+voffcv =0.02
+kt2 = -0.042
+uc1 =0
+jswgs = 1e-010
+bvs = 10
+jswgd = 1e-010
+bvd =10
+mjs = 0.5
+pbswgs = 1
+cjd = 0.0005
+mjswd = 0.33
+tpb = 0.005
+tpbswg =0.005
+toxm = 1.4e-009
+wln = 1
+wwn = 1
+toxref = 1.4e-009
+k3 =0
+dvt1 = 0.52
+dvt2w =0
+dvtp0 = 1e-007
+xj = 2e-008
+phin = 0
+cit =0
+etab = 0
+ub =1.1e-017
+ags = 1e-020
+b1 =0
+pclm =0.18
+drout =0.45
+pscbe2 =1e-007
+pditsl =2.3e+006
+rdw =150
+prwg = 0
+alpha1 =0.005
+cgidl =0.0002
+cigbinv = 0.004
+bigc = 0.0028
+cigsd =0.002
+ntox = 1
+cgdl = 2.495e-10
+acde = 1
+ute =-1.5
+prt =0
+njs = 1
+xjbvs = 1
+njd =1
+xjbvd = 1
+pbsws = 1
+cjswgs = 3e-010
+mjd = 0.5
+pbswgd = 1
+tcj = 0.001
+tcjswg =0.001
+dmcg =0e-006 dmci =0e-006 dmdg = 0e-006 dmcgt = 0e-007
+dwj = 0.0e-008
+rshg = 0.4
+rbps = 15
+xgw = 0e-007
+gbmin = 1e-010
+rbdb = 15
+xgl = 0e-008
+rbpb = 5
+rbsb = 15
+rbpd = 15
+ngcon =1

.MODEL PMOS PMOS LEVEL   = 54
+binunit = 1
+capmod = 2
+diomod = 1
+permod = 1
+tnom = 27
+epsrox = 3.9
+LL =0
+lw =0
+lwl = 0
+vth0 = -0.22
+k3b = 0
+dvt2 = -0.032
+dsub = 0.7
+dvtp1 = 0.05
+ngate =5e+020
+cdsc = 0.000258
+voff =-0.15
+vfb = 0.55
+uc =4.6e-013
+a1 =0
+keta = -0.047
+pdiblc1 = 0.03
+pvag = 1e-020
+fprout =0.2
+rsh = 3
+rdswmin = 0
+prwb = 6.8e-011
+beta0 =30
+egidl = 0.8
+aigbacc = 0.012
+nigbacc = 1
+eigbinv= 1.1
+cigc = 0.0008
+nigc = 1
+xrcrg1 = 12
+cgso = 7.43e-010
+cgsl =1e-014
+moin =15
+kt1 =-0.19
+ua1 =-1e-009
+at = 33000
+paramchk= 1
+igcmod = 1
+rdsmod = 0
+acnqsmod= 0
+toxe = 1.4e-009
+wint = 5e-009
+wl =0
+ww =0
+wwl = 0
+k1 = 0.39
+w0 = 2.5e-006
+dvt0w =0
+minv = 0.05
+lpe0 = 5.75e-008
+ndep =2.8e+018
+cdscb = 0
+nfactor = 2
+u0 = 0.0095
+vsat = 90000
+a2 =1
+dwg =0
+pdiblc2 = 0.0055
+delta =0.014
+pdits =0.2
+rdsw = 250
+rdwmin = 0
+wr =1
+agidl =0.0002
+bigbacc = 0.0028
+aigbinv = 0.014
+nigbinv = 3
+aigsd =0.0087
+poxedge =1
+xrcrg2 = 5
+cgdo =7.43e-010
+ckappas = 0.5
+noff = 0.9
+kt1l =0
+ub1 =2e-018
+mobmod = 0
+igbmod = 1
+rbodymod= 1
+trnqsmod= 0
+toxp =7e-010
+lint = 1.2e-008
+lln =1
+lwn = 1
+xpart =0
+k2 = 0.05
+dvt0 = 3.9
+dvt1w =0
+voffl =0
+lpeb =2.3e-010
+nsd =1e+020
+cdscd =6.1e-008
+eta0 =0.15
+ua = 1.6e-009
+a0 =1.2
+b0 =-1e-020
+dwb =0
+pdiblcb = 3.4e-008
+pscbe1 =8.14e+08
+pditsd =0.23
+rsw = 160
+rswmin = 0
+alpha0 =0.074
+bgidl =2.1e+009
+cigbacc = 0.002
+bigbinv = 0.004
+aigc = 0.69
+bigsd =0.0012
+pigcd = 1
+cgbo =2.56e-011
+ckappad = 0.5
+voffcv =0.02
+kt2 = -0.052
+uc1 =0
+geomod = 1
+rgatemod= 1
+toxm = 1.4e-009
+wln = 1
+wwn = 1
+toxref = 1.4e-009
+k3 =0
+dvt1 = 0.635
+dvt2w =0
+dvtp0 =0.5e-008
+xj = 2e-008
+phin = 0
+cit =0
+etab = 0
+ub = 8e-018
+ags =1e-020
+b1 =0
+pclm = 0.55
+drout =0.56
+pscbe2 =9.58e-07
+pditsl =2.3e+006
+rdw = 160
+prwg = 3.22e-008
+alpha1 =0.005
+cgidl =0.0002
+cigbinv = 0.004
+bigc =0.0012
+cigsd =0.0008
+ntox = 1
+cgdl = 1e-014
+acde = 1
+ute = -1.5
+prt =0
+fnoimod = 1 tnoimod = 0
+jss =0.0001 jsws =1e-011 jswgs = 1e-010 njs =1
+ijthsfwd= 0.01
+jsd = 0.0001
+ijthdfwd= 0.01
+pbs =1
+cjsws =5e-010
+mjswgs =0.33
+pbswd = 1
+cjswgd = 5e-010
+tpbsw =0.005
+xtis = 3
+dmcg = 5e-006
+dwj = 4.5e-008
+rshg = 0.4
+rbps = 15
+ijthsrev= 0.001
+jswd =1e-011
+ijthdrev= 0.001
+cjs = 0.0005
+mjsws = 0.33
+pbd =1
+cjswd =5e-010
+mjswgd = 0.33
+tcjsw =0.001
+xtid = 3
+dmci = 5e-006
+xgw = 3e-007
+gbmin = 1e-010
+rbdb = 15
+bvs =10
+jswgd = 1e-010
+bvd =10
+mjs = 0.5
+pbswgs = 1
+cjd = 0.0005
+mjswd =0.33
+tpb = 0.005
+tpbswg =0.005
+dmdg = 5e-006
+xgl = 4e-008
+rbpb = 5
+rbsb =15
+xjbvs = 1
+njd =1
+xjbvd = 1
+pbsws = 1
+cjswgs = 3e-010
+mjd = 0.5
+pbswgd = 1
+tcj = 0.001
+tcjswg =0.001
+dmcgt =6e-007
+rbpd = 15
+ngcon =1

.control
set color0 =white
set color1=black
op
show all
*Barrido de frecuencia
ac dec 10 1 1ghz
*Impedancia del espejo de corriente ro AC
plot -v(dcasc)/i(vo)
*Impedancia total que ve la fuente AC con el espejo y la resistencia de 100 en serie
plot -v(vo)/i(vo)

.endc


