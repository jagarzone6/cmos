* Simulación Circuito Amplificador Operacional de dos etapas
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

Vdd_1 Vdd_1 0 DC 2.5 AC 0
Vss_1 Vss_1 0 DC -2.5 AC 0

*Vin2_1 vinM2_1 0 DC 0 AC 0
////////////------////////////////////
*Circuito del amplificador operacional de dos etapas
M1_1 drainM1_1 vout_1 sourceM1_1 Vss_1 nmosG W=8e-06 L=1.6e-06
M2_1 drainM2_1 vinM1_1 sourceM1_1 Vss_1 nmosG W=8e-06 L=1.6e-06

M3_1 drainM1_1 drainM1_1 Vdd_1 Vdd_1 pmosG W=1.76e-05 L=1.6e-06
M4_1 drainM2_1 drainM1_1 Vdd_1 Vdd_1 pmosG W=1.76e-05 L=1.6e-06

M5_1 sourceM1_1 vbiasM5_1 Vss_1 Vss_1 nmosG W=3.2e-06 L=1.6e-06

M6_1 vout_1 drainM2_1 Vdd_1 Vdd_1 pmosG W=0.00015999999999999999 L=1.6e-06

M7_1 vout_1 vbiasM5_1 Vss_1 Vss_1 nmosG W=1.92e-05 L=1.6e-06

Cl_1 vout_1 0 10p
Cc_1 vout_1 drainM2_1 4.2239999999999995e-13
////////////------////////////////////
*Circuito espejo ideal
*Iref Espejo N de 0.00023231999999999997 Amps
Iref_1 0 vbiasM5_1 DC 0.00023231999999999997 AC 0
M8_1 vbiasM5_1 vbiasM5_1 Vss_1 Vss_1 nmosG W=3.2e-06 L=1.6e-06
////////////------////////////////////

*Fuente DC en vinM1_1
Vindc_1 vinM1_1 0 DC 0 AC 0

* Modelos para tecnología 0.8u < L < 200u 10u < W < 10000u  Vdd=2.5V (Allen)
* lambda cambia de acuerdo con la longitud del canal
* nMOS: lambda=0.04 para L=1u y lambda=0.01 para L=2u
* pMOS: lambda=0.05 para L=1u y lambda=0.01 para L=2u

.model nmosG nmos level=2
+ vto = 0.7 kp = 110e-6 gamma = 0.4 phi = 0.7
+ tox = 14e-9 cj = 770e-6 cjsw = 380e-12 mj = 0.5 mjsw = 0.38
+ cgso = 220e-12 cgdo = 220e-12 cgbo = 700e-12
+ lambda = 0.04

.model pmosG pmos level=2
+ vto = -0.7 kp = 50e-6 gamma = 0.57 phi = 0.8
+ tox = 14e-9 cj = 560e-6 cjsw = 350e-12 mj = 0.5 mjsw = 0.35
+ cgso = 220e-12 cgdo = 220e-12 cgbo = 700e-12
+ lambda = 0.05

.control
set temp = 0
set tnom = 0
set color0 =white
set color1=black
op
show all

*Simulacion en DC vin vs vout y I(vdd_1) vs vin, para observar la rampa de operacion del amplificador
dc vindc_1 -4 4 0.0001
plot v(vout_1)
plot i(vss_1)
.endc
