*** SPICE deck for cell Current_mirror_bias{sch} from library Fig-20-25-Sim
*** Created on Mon Oct 03, 2016 12:52:34
*** Last revised on Mon Oct 03, 2016 13:26:20
*** Written on Mon Oct 03, 2016 13:28:31 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd

*** TOP LEVEL CELL: Current_mirror_bias{sch}
Mnmos@0 gnd net@13 net@30 gnd NMOS L=2U W=10U
Mnmos@1 gnd net@13 net@13 gnd NMOS L=2U W=10U
Mnmos@3 net@21 net@30 net@13 gnd NMOS L=1U W=10U
Mnmos@4 net@21 net@13 Iref2 gnd NMOS L=2U W=40U
Mpmos@0 net@30 net@30 vdd vdd PMOS L=100U W=10U
Mpmos@1 net@13 net@21 vdd vdd PMOS L=2U W=30U
Mpmos@2 vdd net@21 net@21 vdd PMOS L=2U W=30U
Rres@0 Iref2 gnd 6.5k
.END
