* Bogotá 5 de octubre de 2016
* Universidad Nacional de Colombia 
* CMOS Analógico
* Simulación circuito figura 20.22 Baker (pg 629)
* Grupo Jorge Garzón, Esteban Iafrancesco

VDD VDD 0 DC 1 AC 0
*Vbiasp G4 0 
*Vbiasn D4 0
*Vreg Vreg 0
M1 D1 D1 VDD VDD pmos W=10 L=20
M2 D1 G2 S2 0 nmos W=10 L=1
M3 G4 D1 G2 0 nmos W=10 L=1
M4 D4 G4 VDD VDD pmos W=100 L=2
M5 D4 D4 0 0 nmos W=50 L=2
M6 G6 G6 VDD VDD pmos W=100 L=2
M7 G6 G7 0 0 nmos W=50 L=2
M8 D8 G6 VDD VDD pmos W=100 L=2
M9 D8 D4 0 0 nmos W=50 L=2
M10 G7 D8 VDD VDD pmos W=100 L=2
M11 G7 G7 S11 0 nmos W=50 L=2
R S11 0 5500
D1 G4 VDD POWERMOD AREA=2 W=6um TEMP=100
D2 D4 0 POWERMOD AREA=2 W=6um TEMP=100
.MODEL POWERMOD NUMD LEVEL=2

.MODEL NMOS NMOS LEVEL = 3 NSUB =1E17
+ TOX =200E-10
+ PHI =0.7 VTO = 0.8
+ UO = 650 ETA = 3.0E-6
+ KP=120E-6 VMAX =1E5
+ RSH = 0 NFS =1E12
+ XJ = 500E-9LD = 100E-9
+ CGDO =200E-12 CGSO =200E-12 PB = 1
+ CJ = 400E-6
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.5 DELTA = 3.0 THETA = 0.1 KAPPA =0.3
+ TPG = 1 CGBO =1E-10 MJ = 0.5
*
.MODEL PMOS PMOS LEVEL = 3 NSUB =1E17
+ TOX =200E-10
+ PHI = 0.7 VTO = -0.9 ETA = 0
+ UO = 250 VMAX =5E4
+ KP = 40E-6
+ RSH = 0 NFS =1E12 LD = 100E-9
+ XJ = 500E-9 CGSO =200E-12
+ CGDO =200E-12
+ CJ = 400E-6 PB=1
+ CJSW =300E-12 MJSW =0.5 GAMMA = 0.6 DELTA =0.1 THETA = 0.1 KAPPA = 1
+ TPG = -1 CGBO =1E-10 MJ = 0.5


.control
op
show all
dc VDD 0 1 0.01
plot v(G4) v(D4) 
.endc
	

