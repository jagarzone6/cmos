* Simulación Circuito De las figura 20,15 CMOS Current Mirror Level 3
* Universidad Nacional de Colombia 2016
* CMOS Analógico
* Grupo Jorge Garzón, Esteban Iafrancesco A

Vdd_1 Vdd_1 0 DC 2.5 AC 0
Vss_1 Vss_1 0 DC -2.5 AC 0

////////////------////////////////////
*Circuito del amplificador operacional de dos etapas

M1_1 drainM1_1 vinM1_1 sourceM1_1 Vss_1 nmoslevel3 W=8u L=1.6u
M2_1 drainM2_1 vinM2_1 sourceM1_1 Vss_1 nmoslevel3 W=8u L=1.6u

M3_1 drainM1_1 drainM1_1 Vdd_1 Vdd_1 pmoslevel3 W=12u L=1.6u
M4_1 drainM2_1 drainM1_1 Vdd_1 Vdd_1 pmoslevel3 W=12u L=1.6u

M5_1 sourceM1_1 vbiasM5_1 Vss_1 Vss_1 nmoslevel3 W=1.6u L=1.6u

M6_1 vout_1 drainM2_1 Vdd_1 Vdd_1 pmoslevel3 W=152u L=1.6u

M7_1 vout_1 vbiasM5_1 Vss_1 Vss_1 nmoslevel3 W=9.6u L=1.6u

Cl_1 vout_1 0 10p
Cc_1 vout_1 drainM2_1 3p

////////////------////////////////////
*Circuito del multiplicador beta



VRLref sourceM2 RLo DC 0 AC 0
VM1ref Vm1 0 DC 0 AC 0

* Modelos para tecnología 0.8u < L < 200u 10u < W < 10000u  Vdd=2.5V (Allen)
* lambda cambia de acuerdo con la longitud del canal
* nMOS: lambda=0.04 para L=1u y lambda=0.01 para L=2u
* pMOS: lambda=0.05 para L=1u y lambda=0.01 para L=2u

.model nmoslevel2 nmos level=2
+ vto = 0.7	kp = 110e-6	gamma = 0.4	phi = 0.7
+ tox = 14e-9	cj = 770e-6	cjsw = 380e-12	mj = 0.5	mjsw = 0.38
+ cgso = 220e-12	cgdo = 220e-12	cgbo = 700e-12
+ lambda = 0.04

.model pmoslevel2 pmos level=2
+ vto = -0.7	kp = 50e-6	gamma = 0.57	phi = 0.8
+ tox = 14e-9	cj = 560e-6	cjsw = 350e-12	mj = 0.5	mjsw = 0.35
+ cgso = 220e-12	cgdo = 220e-12	cgbo = 700e-12
+ lambda = 0.05

.tran .1ms 1m uic
.ic v(gatem1)=0 v(drainm2)=0
.control
set color0 =white
set color1=black
op
show all
dc vdd 0 10 0.01
plot i(vrlref) i(vm1ref)
run
plot i(vrlref)
.endc
